module Inst_Rom(
    input [4:0] pc,
    output [31:0] inst
);
    // Define a ROM array to store the instructions
    wire [31:0] rom [0:31]; 

    // Assign values to the instruction ROM
    assign rom[5'h00] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h01] = 32'b000000_00001_00000_00010_00000_100000;  // ADD $v0, $a0, $a1
    assign rom[5'h02] = 32'b000000_00001_00000_00010_00000_100010;  // SUB $v0, $a0, $a2
    assign rom[5'h03] = 32'b000000_00001_00000_00011_00000_100011;  // SUBU $v1, $a0, $a1
    assign rom[5'h04] = 32'b000000_00010_00001_00000_00000_101010;  // SLT $v0, $a1, $a2
    assign rom[5'h05] = 32'b000000_00010_00001_00000_00000_101011;  // SLTU $v0, $a1, $a2
    assign rom[5'h06] = 32'b001111_00000_00110_0000000000000000;  // LUI $a2, 0x0008
    assign rom[5'h07] = 32'b001000_00110_01110_0000000000000100;  // ADDI $a3, $a2, 4
    assign rom[5'h08] = 32'b100011_00110_01000_0000000000000010;  // LW $t0, 2($a3)
    assign rom[5'h09] = 32'b101011_00000_00010_0000000000000010;  // SW $v0, 2($v0)
    assign rom[5'h0A] = 32'b000100_00001_00000_0000000000000001;  // BEQ $v1, $v0, 1
    assign rom[5'h0B] = 32'b000100_00001_00000_0000000000000001;  // BEQ $v1, $a0, 1
    assign rom[5'h0C] = 32'b000010_00000000000000000000001000;  // J 0x00000008
    assign rom[5'h0D] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h0E] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h0F] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h10] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h11] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h12] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h13] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h14] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h15] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h16] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h17] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h18] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h19] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h1A] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h1B] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h1C] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h1D] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h1E] = 32'b000000_00000_00000_00000_00000_000000;  // NOP
    assign rom[5'h1F] = 32'b000000_00000_00000_00000_00000_000000;  // NOP

    // Output the instruction based on the pc (program counter)
    assign inst = rom[pc];

endmodule
